// Vendor 		: 
// Author 		: ling
// Filename 	: bus_checker 
// Date Created: 2022.04.26 
// Version		: V1.0
// File description	:
// Revision History :

`include "axi_base_base_vseq.sv"
`include "axi_base_random_vseq.sv"
`include "axi_base_random_reset_vseq.sv"
`include "axi_base_disabled_vseq.sv"
`include "axi_base_cfg_update_on_fly_vseq.sv"
`include "axi_base_common_vseq.sv"
`include "axi_base_stress_all_vseq.sv"
