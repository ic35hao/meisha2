// *************************************************************************************************
// Vendor 		: 
// Author 		: ling
// Filename 	: mst_port_info 
// Date Created: 2022.05.01 
// Version		: V1.0
// -------------------------------------------------------------------------------------------------
// File description	:
// -------------------------------------------------------------------------------------------------
// Revision History :
// *************************************************************************************************

//--------------------------------------------------------------------------------------------------
// module declaration
//--------------------------------------------------------------------------------------------------

class mst_port_info extends bind_abs_pkg::base_port_info;

    access_addr_info acc_info;
    //----------------------------------------------------------------------------------------------
    // Parameter Define
    //----------------------------------------------------------------------------------------------
    `uvm_object_utils(mst_port_info)
    


// Constructor: new
extern function new(string name = "mst_port_info");

endclass: mst_port_info

function mst_port_info::new(string name = "mst_port_info");
    super.new(name);
endfunction: new
//--------------------------------------------------------------------------------------------------
// eof
//--------------------------------------------------------------------------------------------------