// *************************************************************************************************
// Vendor 		: 
// Author 		: ling
// Filename 	: apb_port_info 
// Date Created: 2022.04.27 
// Version		: V1.0
// -------------------------------------------------------------------------------------------------
// File description	:
// -------------------------------------------------------------------------------------------------
// Revision History :
// *************************************************************************************************

//--------------------------------------------------------------------------------------------------
// module declaration
//--------------------------------------------------------------------------------------------------

class apb_port_info extends base_port_info;

    //----------------------------------------------------------------------------------------------
    // Parameter Define
    //----------------------------------------------------------------------------------------------
    //`uvm_object_utils(apb_port_info)

    `uvm_object_new

endclass: apb_port_info
