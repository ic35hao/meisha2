// *************************************************************************************************
// Vendor 		: 
// Author 		: ling
// Filename 	: axi_port_info 
// Date Created: 2022.04.27 
// Version		: V1.0
// -------------------------------------------------------------------------------------------------
// File description	:
// -------------------------------------------------------------------------------------------------
// Revision History :
// *************************************************************************************************

//--------------------------------------------------------------------------------------------------
// module declaration
//--------------------------------------------------------------------------------------------------

class axi_port_info extends base_port_info;

    //----------------------------------------------------------------------------------------------
    // Parameter Define
    //----------------------------------------------------------------------------------------------
    //`uvm_object_utils(axi_port_info)

    `uvm_object_new

endclass: axi_port_info