

class tlul_base_virtual_sequencer extends cip_base_virtual_sequencer #(.CFG_T(tlul_base_env_cfg), .COV_T(tlul_base_env_cov));
  `uvm_component_utils(tlul_base_virtual_sequencer)

  `uvm_component_new

endclass
